// Copyright (C) 2016  Intel Corporation. All rights reserved.
//
// Your use of Intel Corporation's design tools, logic functions and
// other software and tools, and its AMPP partner logic functions, and
// any output files from any of the foregoing (including device
// programming or simulation files), and any associated documentation
// or information are expressly subject to the terms and conditions of
// the Intel Program License Subscription Agreement, the Intel Quartus
// Prime License Agreement, the Intel MegaCore Function License
// Agreement, or other applicable license agreement, including,
// without limitation, that your use is for the sole purpose of
// programming logic devices manufactured by Intel and sold by Intel
// or its authorized distributors.  Please refer to the applicable
// agreement for further details.

// Generated by Quartus.
// With edits from Matthew Naylor, August 2019.

// True dual-port block RAM
// ========================

module BlockRAMTrueDualMixed (
  ADDR_A,
  ADDR_B,
  CLK,
  DI_A,
  DI_B,
  WE_A,
  WE_B,
  DO_A,
  DO_B
  );

  parameter ADDR_WIDTH_A = 1;
  parameter ADDR_WIDTH_B = 1;
  parameter DATA_WIDTH_A = 1;
  parameter NUM_ELEMS    = 1;
  parameter RD_DURING_WR = "OLD_DATA";     // Or: "DONT_CARE"
  parameter DO_REG_A     = "UNREGISTERED"; // Or: "CLOCK0"
  parameter DO_REG_B     = "UNREGISTERED"; // Or: "CLOCK0"
  parameter INIT_FILE    = "UNUSED";
  parameter DEV_FAMILY   = "Stratix V";

  localparam RATIO = 1 << (ADDR_WIDTH_A - ADDR_WIDTH_B);
  localparam DATA_WIDTH_B = DATA_WIDTH_A * RATIO;

  input [ADDR_WIDTH_A-1:0] ADDR_A;
  input [ADDR_WIDTH_B-1:0] ADDR_B;
  input CLK;
  input [DATA_WIDTH_A-1:0] DI_A;
  input [DATA_WIDTH_B-1:0] DI_B;
  input WE_A;
  input WE_B;
  output [15:0] DO_A;
  output [7:0] DO_B;

  altsyncram  altsyncram_component (
        .address_a (ADDR_A),
        .address_b (ADDR_B),
        .clock0 (CLK),
        .data_a (DI_A),
        .data_b (DI_B),
        .wren_a (WE_A),
        .wren_b (WE_B),
        .q_a (DO_A),
        .q_b (DO_B),
        .aclr0 (1'b0),
        .aclr1 (1'b0),
        .addressstall_a (1'b0),
        .addressstall_b (1'b0),
        .byteena_a (1'b1),
        .byteena_b (1'b1),
        .clock1 (1'b1),
        .clocken0 (1'b1),
        .clocken1 (1'b1),
        .clocken2 (1'b1),
        .clocken3 (1'b1),
        .eccstatus (),
        .rden_a (1'b1),
        .rden_b (1'b1));
  defparam
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.intended_device_family = DEV_FAMILY,
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.numwords_a = 2**ADDR_WIDTH_A,
    altsyncram_component.numwords_b = 2**ADDR_WIDTH_B,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_a = DO_REG_A,
    altsyncram_component.outdata_reg_b = DO_REG_B,
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.read_during_write_mode_mixed_ports = RD_DURING_WR,
    altsyncram_component.read_during_write_mode_port_a = "NEW_DATA_NO_NBE_READ",
    altsyncram_component.read_during_write_mode_port_b = "NEW_DATA_NO_NBE_READ",
    altsyncram_component.widthad_a = ADDR_WIDTH_A,
    altsyncram_component.widthad_b = ADDR_WIDTH_B,
    altsyncram_component.width_a = DATA_WIDTH_A,
    altsyncram_component.width_b = DATA_WIDTH_B,
    altsyncram_component.width_byteena_a = 1,
    altsyncram_component.width_byteena_b = 1,
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0";

endmodule
